LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY notnbit IS
	GENERIC(
		n : IN NATURAL := 16
	);

	PORT(
		a : IN STD_LOGIC_VECTOR(n-1 DOWNTO 0);
		q : OUT STD_LOGIC_VECTOR(n-1 DOWNTO 0)
	);
END;

ARCHITECTURE bhv OF notnbit IS
BEGIN

	PROCESS
	BEGIN
		nottobe : FOR i IN 0 TO n-1 LOOP
			q(i) <= (NOT a(i));
		END LOOP;
	END PROCESS;

END;
