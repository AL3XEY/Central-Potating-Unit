﻿LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY reg1bit IS
	PORT(
		d, clk : IN STD_LOGIC;
		q : OUT STD_LOGIC
	);
END;

ARCHITECTURE dlatch OF reg1bit IS
BEGIN

END;