LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY cpu16bits IS
	PORT(
		run, resetn, clk : IN STD_LOGIC;
		din : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		busio : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		done : OUT STD_LOGIC
	);
END;

ARCHITECTURE bhv OF cpu16bits IS
BEGIN

END;